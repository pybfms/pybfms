/****************************************************************************
 * simple_bfm_top.sv
 ****************************************************************************/
 
/**
 * Module: simple_bfm_top
 * 
 * TODO: Add module documentation
 */
module simple_bfm_top(input clk);
	
	initial begin
		$display("Hello World");
	end

	simple_bfm bfm_0 (clk);


endmodule


