/****************************************************************************
 * ${bfm}_api_pkg.sv
 ****************************************************************************/
package ${bfm}_api_pkg;
	
	class ${bfm}_api;
${bfm_class_api}
	endclass
	
endpackage
